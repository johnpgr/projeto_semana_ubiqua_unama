module main


pub struct User {
pub mut:
	name string
	email string
	hashed_password string
}
